.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C1608C0G2A100D080AA_p.mod"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/FMMT597.spice.txt"
.include "models/SMAZ15.spice.txt"
.include "models/ZXCT1008F.spice.txt"
XU3 /PWR_IN /SN C1608C0G2A100D080AA_p
R3 /PWR_IN /PWR_OUT {RSENSE1}
R4 /PWR_IN /PWR_OUT {RSENSE2}
XU2 /SN /PWR_IN /COCM ZXCT1008F
R7 /PWR_OUT /SN {RLIM}
I1 /PWR_OUT 0 {ILOAD}
V1 /PWR_IN 0 {VSOURCE}
Q1 /FILTER /BASE /COCM FMMT597
XU1 /BASE /PWR_IN SMAZ15
R5 /FILTER 0 {RSET1}
R6 /FILTER 0 {RSET2}
R1 /BASE 0 {RBASE}
R2 /OUT /FILTER {RFILTER}
XU4 0 /OUT DI_BZX84C4V7
XU5 /OUT 0 C2012C0G2A102J060AA_p
.end
