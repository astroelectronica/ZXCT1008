.title KiCad schematic
.include "C:/AE/ZXCT1008/_models/BZX84C4V7.spice.txt"
.include "C:/AE/ZXCT1008/_models/C1608C0G2A100D080AA_p.mod"
.include "C:/AE/ZXCT1008/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1008/_models/FMMT597.spice.txt"
.include "C:/AE/ZXCT1008/_models/SMAZ15.spice.txt"
.include "C:/AE/ZXCT1008/_models/ZXCT1008F.spice.txt"
R7 /PWR_OUT /SN {RLIM}
I1 /PWR_OUT 0 {ILOAD}
XU1 /BASE /PWR_IN SMAZ15
XU3 /PWR_IN /SN C1608C0G2A100D080AA_p
Q1 /FILTER /BASE /COCM FMMT597
XU2 /SN /PWR_IN /COCM ZXCT1008F
R5 /FILTER 0 {RSET1}
R6 /FILTER 0 {RSET2}
R4 /PWR_IN /PWR_OUT {RSENSE2}
R3 /PWR_IN /PWR_OUT {RSENSE1}
V1 /PWR_IN 0 {VSOURCE}
R1 /BASE 0 {RBASE}
R2 /OUT /FILTER {RFILTER}
XU4 0 /OUT DI_BZX84C4V7
XU5 /OUT 0 C2012C0G2A102J060AA_p
.end
